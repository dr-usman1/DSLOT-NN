module And_Mult_Array(
  input reg [15:0] activation_0, input reg weight_0,
  input reg [15:0] activation_1, input reg weight_1,
  input reg [15:0] activation_2, input reg weight_2,
  input reg [15:0] activation_3, input reg weight_3,
  input reg [15:0] activation_4, input reg weight_4,
  input reg [15:0] activation_5, input reg weight_5,
  input reg [15:0] activation_6, input reg weight_6,
  input reg [15:0] activation_7, input reg weight_7,
  input reg [15:0] activation_8, input reg weight_8,
  input reg [15:0] activation_9, input reg weight_9,
  input reg [15:0] activation_10, input reg weight_10,
  input reg [15:0] activation_11, input reg weight_11,
  input reg [15:0] activation_12, input reg weight_12,
  input reg [15:0] activation_13, input reg weight_13,
  input reg [15:0] activation_14, input reg weight_14,
  input reg [15:0] activation_15, input reg weight_15,
  input reg [15:0] activation_16, input reg weight_16,
  input reg [15:0] activation_17, input reg weight_17,
  input reg [15:0] activation_18, input reg weight_18,
  input reg [15:0] activation_19, input reg weight_19,
  input reg [15:0] activation_20, input reg weight_20,
  input reg [15:0] activation_21, input reg weight_21,
  input reg [15:0] activation_22, input reg weight_22,
  input reg [15:0] activation_23, input reg weight_23,
  input reg [15:0] activation_24, input reg weight_24,
  input reg [15:0] activation_25, input reg weight_25,
  input reg [15:0] activation_26, input reg weight_26,
  input reg [15:0] activation_27, input reg weight_27,
  input reg [15:0] activation_28, input reg weight_28,
  input reg [15:0] activation_29, input reg weight_29,
  input reg [15:0] activation_30, input reg weight_30,
  input reg [15:0] activation_31, input reg weight_31,
  output  [15:0] result_0,  result_1,
  output  [15:0] result_2,  result_3,
  output  [15:0] result_4,  result_5,
  output  [15:0] result_6,  result_7,
  output  [15:0] result_8,  result_9,
  output  [15:0] result_10, result_11,
  output  [15:0] result_12, result_13,
  output  [15:0] result_14, result_15,
  output  [15:0] result_16, result_17,
  output  [15:0] result_18, result_19,
  output  [15:0] result_20, result_21,
  output  [15:0] result_22, result_23,
  output  [15:0] result_24, result_25,
  output  [15:0] result_26, result_27,
  output  [15:0] result_28, result_29,
  output  [15:0] result_30, result_31
);

  ActivationMultiplier inst_0 (
    .activation(activation_0),
    .weight(weight_0),
    .result(result_0)
  );
  
  ActivationMultiplier inst_1 (
    .activation(activation_1),
    .weight(weight_1),
    .result(result_1)
  );

ActivationMultiplier inst_2 (
.activation(activation_2),
.weight(weight_2),
.result(result_2)
);

ActivationMultiplier inst_3 (
.activation(activation_3),
.weight(weight_3),
.result(result_3)
);

ActivationMultiplier inst_4 (
.activation(activation_4),
.weight(weight_4),
.result(result_4)
);

ActivationMultiplier inst_5 (
.activation(activation_5),
.weight(weight_5),
.result(result_5)
);

ActivationMultiplier inst_6 (
.activation(activation_6),
.weight(weight_6),
.result(result_6)
);

ActivationMultiplier inst_7 (
.activation(activation_7),
.weight(weight_7),
.result(result_7)
);

ActivationMultiplier inst_8 (
.activation(activation_8),
.weight(weight_8),
.result(result_8)
);

ActivationMultiplier inst_9 (
.activation(activation_9),
.weight(weight_9),
.result(result_9)
);

ActivationMultiplier inst_10 (
.activation(activation_10),
.weight(weight_10),
.result(result_10)
);

ActivationMultiplier inst_11 (
.activation(activation_11),
.weight(weight_11),
.result(result_11)
);

ActivationMultiplier inst_12 (
.activation(activation_12),
.weight(weight_12),
.result(result_12)
);

ActivationMultiplier inst_13 (
.activation(activation_13),
.weight(weight_13),
.result(result_13)
);

ActivationMultiplier inst_14 (
.activation(activation_14),
.weight(weight_14),
.result(result_14)
);

ActivationMultiplier inst_15 (
.activation(activation_15),
.weight(weight_15),
.result(result_15)
);

ActivationMultiplier inst_16 (
.activation(activation_16),
.weight(weight_16),
.result(result_16)
);

ActivationMultiplier inst_17 (
.activation(activation_17),
.weight(weight_17),
.result(result_17)
);

ActivationMultiplier inst_18 (
.activation(activation_18),
.weight(weight_18),
.result(result_18)
);

ActivationMultiplier inst_19 (
.activation(activation_19),
.weight(weight_19),
.result(result_19)
);

ActivationMultiplier inst_20 (
.activation(activation_20),
.weight(weight_20),
.result(result_20)
);

ActivationMultiplier inst_21 (
.activation(activation_21),
.weight(weight_21),
.result(result_21)
);

ActivationMultiplier inst_22 (
.activation(activation_22),
.weight(weight_22),
.result(result_22)
);

ActivationMultiplier inst_23 (
.activation(activation_23),
.weight(weight_23),
.result(result_23)
);

ActivationMultiplier inst_24 (
.activation(activation_24),
.weight(weight_24),
.result(result_24)
);

ActivationMultiplier inst_25 (
.activation(activation_25),
.weight(weight_25),
.result(result_25)
);

ActivationMultiplier inst_26 (
.activation(activation_26),
.weight(weight_26),
.result(result_26)
);

ActivationMultiplier inst_27 (
.activation(activation_27),
.weight(weight_27),
.result(result_27)
);

ActivationMultiplier inst_28 (
.activation(activation_28),
.weight(weight_28),
.result(result_28)
);

ActivationMultiplier inst_29 (
.activation(activation_29),
.weight(weight_29),
.result(result_29)
);

ActivationMultiplier inst_30 (
.activation(activation_30),
.weight(weight_30),
.result(result_30)
);

ActivationMultiplier inst_31 (
.activation(activation_31),
.weight(weight_31),
.result(result_31)
);

endmodule
